`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    14:36:52 09/30/2016 
// Design Name: 
// Module Name:    RippleCarryAdder 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module RippleCarryAdder(a, b, cin, sum, cout);

input [15:0] a;
input [15:0] b;
input cin;

output [15:0]sum;
output cout;

wire[14:0] c;

FullAdder a1(a[0],b[0],cin,sum[0],c[0]);
FullAdder a2(a[1],b[1],c[0],sum[1],c[1]);
FullAdder a3(a[2],b[2],c[1],sum[2],c[2]);
FullAdder a4(a[3],b[3],c[2],sum[3],c[3]);
FullAdder a5(a[4],b[4],c[3],sum[4],c[4]);
FullAdder a6(a[5],b[5],c[4],sum[5],c[5]);
FullAdder a7(a[6],b[6],c[5],sum[6],c[6]);
FullAdder a8(a[7],b[7],c[6],sum[7],c[7]);
FullAdder a9(a[8],b[8],c[7],sum[8],c[8]);
FullAdder a10(a[9],b[9],c[8],sum[9],c[9]);
FullAdder a11(a[10],b[10],c[9],sum[10],c[10]);
FullAdder a12(a[11],b[11],c[10],sum[11],c[11]);
FullAdder a13(a[12],b[12],c[11],sum[12],c[12]);
FullAdder a14(a[13],b[13],c[12],sum[13],c[13]);
FullAdder a15(a[14],b[14],c[13],sum[14],c[14]);
FullAdder a16(a[15],b[15],c[14],sum[15],cout);

endmodule